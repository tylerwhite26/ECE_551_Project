module ble_module()
    // Placeholder for BLE module
    // Should send 'G' and 'S' to AUTH_blk to turn the segway on and off.
    // 'G' asserts PWR_UP and 'S' deasserts PWR_UP when rider_off is high.
    
endmodule